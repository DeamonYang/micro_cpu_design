`timaecale 1ns/1ps
/****************************************************************
@file name	: mem_stage.sv
@description: mem  control top wrapper
=================================================================
revision		data		author		commit
  0.1		2019/11/16	  deamonyang	draft
****************************************************************/